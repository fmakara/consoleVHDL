library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
entity ROM_DESSINS is Port (
	CLK      : in  STD_LOGIC;
	RESET    : in  STD_LOGIC;
	ADDR_OUT : in  STD_LOGIC_VECTOR (9 downto 0);
	DATA_OUT : out STD_LOGIC_VECTOR (17 downto 0);
	ADDR_IN  : in  STD_LOGIC_VECTOR (9 downto 0);
	DATA_IN  : in STD_LOGIC_VECTOR (17 downto 0);
	WE       : in  STD_LOGIC
); 
end ROM_DESSINS;
architecture Behavioral of ROM_DESSINS is
TYPE memoire IS ARRAY(0 to 1023) OF STD_LOGIC_VECTOR(17 downto 0);--RAMBLOCK 
SIGNAL M : memoire := (
	"000100001111110000","000010101111100110","000011101111011000","000011101111001010",
	"000011101110111100","000100011110101011","000100011110011010","000010111110001111",
	"000100011101111110","000100011101101101","000001011101101000","011111001011101100",
	"011111001001110000","011111000111110100","001011100111000110","100101100100110000",
	"001000110100001101","010011010011000000","011010010001010111","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","111000000000000000",
	"111000000100000000","111000001000000000","111000001100000000","111000010000000000",
	"111000010100000000","111000011000000000","111000011100000000","111000100000000000",
	"111000100100000000","111000101000000000","111000101100000000","111000110000000000",
	"111000110100000000","111000111000000000","111000111100000000","111001000000000000",
	"111001000100000000","111001001000000000","111001001100000000","111001010000000000",
	"111001010100000000","111001011000000000","111001011100000000","111001100000000000",
	"111001100100000000","111001101000000000","111001101100000000","111001110000000000",
	"111001110100000000","111001111000000000","111001111100000000","111010000000000000",
	"111010000100000000","111010001000000000","111010001100000000","111010010000000000",
	"111010010100000000","111010011000000000","111010011100000000","111010100000000000",
	"111010100100000000","111010101000000000","111010101100000000","111010110000000000",
	"111010110100000000","111010111000000000","111010111100000000","111011000000000000",
	"111011000100000000","111011001000000000","111011001100000000","111011010000000000",
	"111011010100000000","111011011000000000","111011011100000000","111011100000000000",
	"111011100100000000","111011101000000000","111011101100000000","111011110000000000",
	"111011110100000000","111011111000000000","111011111100000000","111100000000000000",
	"111100000100000000","111100001000000000","111100001100000000","111100010000000000",
	"111100010100000000","111100011000000000","111100011100000000","111100100000000000",
	"111100100100000000","111100101000000000","111100101100000000","111100110000000000",
	"111100110100000000","111100111000000000","111100111100000000","111101000000000000",
	"111101000100000000","111101001000000000","111101001100000000","111101010000000000",
	"111101010100000000","111101011000000000","111101011100000000","111101100000000000",
	"111101100100000000","111101101000000000","111101101100000000","111101110000000000",
	"111101110100000000","111101111000000000","111101111100000000","111110000000000000",
	"111110000100000000","111110001000000000","111110001100000000","111110010000000000",
	"111110010100000000","111110011000000000","111110011100000000","111110100000000000",
	"111000001000000000","111000000100000001","111000001000000001","111000000100000010",
	"111000001000000010","111000000100000011","111000001000000011","111000000000000100",
	"111000000100000100","111000001000000100","111000000000000101","111000000100000101",
	"111000001000000101","111000000000000110","111000000100000110","111000001000000110",
	"111000000000000111","111000000100000111","111000001000000111","111000000000001000",
	"111000000100001000","111000001000001000","111000000000001001","111000000100001001",
	"111000001000001001","111000000000001010","111000000100001010","111000001000001010",
	"111000000000001011","111000000100001011","111000001000001011","111000000000001100",
	"111000000100001100","111000001000001100","111000000000001101","111000000100001101",
	"111000001000001101","111000000000001110","111000000100001110","111000001000001110",
	"111000000000001111","111000000100001111","111000001000001111","111000000000010000",
	"111000000100010000","111000001000010000","111000000000010001","111000000100010001",
	"111000001000010001","111000000000010010","111000000100010010","111000001000010010",
	"111000000000010011","111000000100010011","111000001000010011","111000000000010100",
	"111000000100010100","111000001000010100","111000000000010101","111000000100010101",
	"111000001000010101","111000000000010110","111000000100010110","111000001000010110",
	"111000000000010111","111000000100010111","111000001000010111","111000000000011000",
	"111000000100011000","111000001000011000","111000000100011001","111000001000011001",
	"111000000100011010","111000001000011010","111000000100011011","111000001000011011",
	"111000001000011100","001000000000000000","001000000100000000","001000001000000000",
	"001000001100000000","001000010000000000","001000010100000000","001000011000000000",
	"001000011000000001","001000011000000010","001000011000000011","001000011000000100",
	"001000000000000101","001000000100000101","001000001000000110","001000001100000110",
	"001000010000000111","001000010100000111","001000011000001000","001000010000001001",
	"001000010100001001","001000001000001010","001000001100001010","001000000000001011",
	"001000000100001011","001000000000001101","001000000100001101","001000001000001101",
	"001000001100001101","001000010000001101","001000010100001101","001000011000001101",
	"001000011000001110","001000011000001111","001000011000010000","001000011000010001",
	"111000000000000000","111000000000000001","111000000000000010","111000000000000011",
	"111000000000000100","111000000000000101","111000000000000110","111000000000000111",
	"111000000000001000","111000000000001001","111000000000001010","111000000000001011",
	"111000000000001100","111000000000001101","111000000000001110","111000000000001111",
	"111000000000010000","111000000000010001","111000000000010010","111000000000010011",
	"111000000000010100","111000000000010101","111000000000010110","111000000000010111",
	"111000000000011000","111000000000011001","111000000000011010","111000000000011011",
	"111000000000011100","111000000000011101","111000000000011110","111000000000011111",
	"111000000000100000","111000000000100001","111000000000100010","111000000000100011",
	"111000000000100100","111000000000100101","111000000000100110","111000000000100111",
	"111000000000101000","111000000000101001","111000000000101010","111000000000101011",
	"111000000000101100","111000000000101101","111000000000101110","111000000000101111",
	"111000000000110000","111000000000110001","111000000000110010","111000000000110011",
	"111000000000110100","111000000000110101","111000000000110110","111000000000110111",
	"111000000000111000","111000000000111001","111000000000111010","111000000000111011",
	"111000000000111100","111000000000111101","111000000000111110","111000000000111111",
	"111000000001000000","111000000001000001","111000000001000010","111000000001000011",
	"111000000001000100","111000000001000101","111000000001000110","111000000001000111",
	"111000000001001000","111000000001001001","111000000001001010","111000000001001011",
	"111000000001001100","111000000001001101","111000000001001110","111000000001001111",
	"111000000001010000","111000000001010001","111000000001010010","111000000001010011",
	"111000000001010100","111000000001010101","111000000001010110","111000000001010111",
	"111000000001011000","111000000001011001","111000000001011010","111000000001011011",
	"111000000001011100","111000000001011101","111000000001011110","111000000001011111",
	"111000000001100000","111000000001100001","111000000001100010","111000000001100011",
	"111000000001100100","111000000001100101","111000000001100110","111000000001100111",
	"111000000001101000","111000000001101001","111000000001101010","111000000001101011",
	"111000000001101100","111000000001101101","111000000001101110","111000000001101111",
	"111000000001110000","111000000001110001","111000000001110010","111000000001110011",
	"111000000001110100","111000000001110101","111000000001110110","111000000001110111",
	"111000000001111000","111000000001111001","111000000001111010","111000000001111011",
	"111000000001111100","111000000001111101","111000000001111110","111000000001111111",
	"111000000010000000","111000000010000001","111000000010000010","111000000010000011",
	"111000000010000100","111000000010000101","111000000010000110","111000000010000111",
	"111000000010001000","111000000010001001","111000000010001010","111000000010001011",
	"111000000010001100","111000000010001101","111000000010001110","111000000010001111",
	"111000000010010000","111000000010010001","111000000010010010","111000000010010011",
	"111000000010010100","111000000010010101","100000000100000000","100000001000000000",
	"100000001100000000","100000000000000001","100000000100000001","100000001000000001",
	"100000001100000001","100000010000000001","100000000000000010","100000000100000010",
	"100000001000000010","100000001100000010","100000010000000010","100000010100000010",
	"100000000100000011","100000001000000011","100000001100000011","100000010000000011",
	"100000010100000011","100000011000000011","100000001000000100","100000001100000100",
	"100000010000000100","100000010100000100","100000011000000100","100000011100000100",
	"100000000100000101","100000001000000101","100000001100000101","100000010000000101",
	"100000010100000101","100000011000000101","100000000000000110","100000000100000110",
	"100000001000000110","100000001100000110","100000010000000110","100000010100000110",
	"100000000000000111","100000000100000111","100000001000000111","100000001100000111",
	"100000010000000111","100000000100001000","100000001000001000","100000001100001000",
	"100000000100000000","100000001000000000","100000001100000000","100000010000000000",
	"100000010100000000","100000011000000000","100000000000000001","101000000100000001",
	"101000001000000001","101000001100000001","101000010000000001","101000010100000001",
	"101000011000000001","100000011100000001","100000000000000010","101000000100000010",
	"101000001000000010","101000001100000010","101000010000000010","101000010100000010",
	"101000011000000010","100000011100000010","100000000000000011","101000000100000011",
	"101000001000000011","101000001100000011","101000010000000011","101000010100000011",
	"101000011000000011","100000011100000011","100000000000000100","101000000100000100",
	"101000001000000100","101000001100000100","101000010000000100","101000010100000100",
	"101000011000000100","100000011100000100","100000000000000101","101000000100000101",
	"101000001000000101","101000001100000101","101000010000000101","101000010100000101",
	"101000011000000101","100000011100000101","100000000000000110","101000000100000110",
	"101000001000000110","101000001100000110","101000010000000110","101000010100000110",
	"101000011000000110","100000011100000110","100000000000000111","101000000100000111",
	"101000001000000111","101000001100000111","101000010000000111","101000010100000111",
	"101000011000000111","100000011100000111","100000000000001000","101000000100001000",
	"101000001000001000","101000001100001000","101000010000001000","101000010100001000",
	"101000011000001000","100000011100001000","100000000000001001","101000000100001001",
	"101000001000001001","101000001100001001","101000010000001001","101000010100001001",
	"101000011000001001","100000011100001001","100000000000001010","101000000100001010",
	"101000001000001010","101000001100001010","101000010000001010","101000010100001010",
	"101000011000001010","100000011100001010","100000000000001011","101000000100001011",
	"101000001000001011","101000001100001011","101000010000001011","101000010100001011",
	"101000011000001011","100000011100001011","100000000000001100","101000000100001100",
	"101000001000001100","101000001100001100","101000010000001100","101000010100001100",
	"101000011000001100","100000011100001100","100000000000001101","101000000100001101",
	"101000001000001101","101000001100001101","101000010000001101","101000010100001101",
	"101000011000001101","100000011100001101","100000000000001110","101000000100001110",
	"101000001000001110","101000001100001110","101000010000001110","101000010100001110",
	"101000011000001110","100000011100001110","100000000100001111","100000001000001111",
	"100000001100001111","100000010000001111","100000010100001111","100000011000001111",
	"001000000100000000","001000001000000000","001000001100000000","001000010000000000",
	"001000010100000000","001000011000000000","001000000000000001","011000000100000001",
	"011000001000000001","011000001100000001","011000010000000001","011000010100000001",
	"011000011000000001","001000011100000001","001000000000000010","011000000100000010",
	"011000001000000010","011000001100000010","011000010000000010","011000010100000010",
	"011000011000000010","001000011100000010","001000000000000011","011000000100000011",
	"011000001000000011","011000001100000011","011000010000000011","011000010100000011",
	"011000011000000011","001000011100000011","001000000000000100","011000000100000100",
	"011000001000000100","011000001100000100","011000010000000100","011000010100000100",
	"011000011000000100","001000011100000100","001000000000000101","011000000100000101",
	"011000001000000101","011000001100000101","011000010000000101","011000010100000101",
	"011000011000000101","001000011100000101","001000000000000110","011000000100000110",
	"011000001000000110","011000001100000110","011000010000000110","011000010100000110",
	"011000011000000110","001000011100000110","001000000000000111","011000000100000111",
	"011000001000000111","011000001100000111","011000010000000111","011000010100000111",
	"011000011000000111","001000011100000111","001000000000001000","011000000100001000",
	"011000001000001000","011000001100001000","011000010000001000","011000010100001000",
	"011000011000001000","001000011100001000","001000000000001001","011000000100001001",
	"011000001000001001","011000001100001001","011000010000001001","011000010100001001",
	"011000011000001001","001000011100001001","001000000000001010","011000000100001010",
	"011000001000001010","011000001100001010","011000010000001010","011000010100001010",
	"011000011000001010","001000011100001010","001000000000001011","011000000100001011",
	"011000001000001011","011000001100001011","011000010000001011","011000010100001011",
	"011000011000001011","001000011100001011","001000000000001100","011000000100001100",
	"011000001000001100","011000001100001100","011000010000001100","011000010100001100",
	"011000011000001100","001000011100001100","001000000000001101","011000000100001101",
	"011000001000001101","011000001100001101","011000010000001101","011000010100001101",
	"011000011000001101","001000011100001101","001000000000001110","011000000100001110",
	"011000001000001110","011000001100001110","011000010000001110","011000010100001110",
	"011000011000001110","001000011100001110","001000000100001111","001000001000001111",
	"001000001100001111","001000010000001111","001000010100001111","001000011000001111",
	"110000000100000000","110000001000000000","110000001100000000","110000010000000000",
	"110000010100000000","110000011000000000","110000000000000001","010000000100000001",
	"010000001000000001","010000001100000001","010000010000000001","010000010100000001",
	"010000011000000001","110000011100000001","110000000000000010","010000000100000010",
	"010000001000000010","010000001100000010","010000010000000010","010000010100000010",
	"010000011000000010","110000011100000010","110000000000000011","010000000100000011",
	"010000001000000011","010000001100000011","010000010000000011","010000010100000011",
	"010000011000000011","110000011100000011","110000000000000100","010000000100000100",
	"010000001000000100","010000001100000100","010000010000000100","010000010100000100",
	"010000011000000100","110000011100000100","110000000000000101","010000000100000101",
	"010000001000000101","010000001100000101","010000010000000101","010000010100000101",
	"010000011000000101","110000011100000101","110000000000000110","010000000100000110",
	"010000001000000110","010000001100000110","010000010000000110","010000010100000110",
	"010000011000000110","110000011100000110","110000000000000111","010000000100000111",
	"010000001000000111","010000001100000111","010000010000000111","010000010100000111",
	"010000011000000111","110000011100000111","110000000000001000","010000000100001000",
	"010000001000001000","010000001100001000","010000010000001000","010000010100001000",
	"010000011000001000","110000011100001000","110000000000001001","010000000100001001",
	"010000001000001001","010000001100001001","010000010000001001","010000010100001001",
	"010000011000001001","110000011100001001","110000000000001010","010000000100001010",
	"010000001000001010","010000001100001010","010000010000001010","010000010100001010",
	"010000011000001010","110000011100001010","110000000000001011","010000000100001011",
	"010000001000001011","010000001100001011","010000010000001011","010000010100001011",
	"010000011000001011","110000011100001011","110000000000001100","010000000100001100",
	"010000001000001100","010000001100001100","010000010000001100","010000010100001100",
	"010000011000001100","110000011100001100","110000000000001101","010000000100001101",
	"010000001000001101","010000001100001101","010000010000001101","010000010100001101",
	"010000011000001101","110000011100001101","110000000000001110","010000000100001110",
	"010000001000001110","010000001100001110","010000010000001110","010000010100001110",
	"010000011000001110","110000011100001110","110000000100001111","110000001000001111",
	"110000001100001111","110000010000001111","110000010100001111","110000011000001111",
	"111000000100000000","111000000000000001","111000000100000001","111000001000000001",
	"111000000100000010","110000000100000000","110000001000000000","110000010100000000",
	"110000000000000001","110000001100000001","110000011000000001","110000000000000010",
	"110000001100000010","110000011000000010","110000000000000011","110000001100000011",
	"110000011000000011","110000000100000100","110000001000000100","110000001100000100",
	"110000010000000100","110000010100000100","110000000100000000","110000001000000000",
	"110000010000000000","110000010100000000","110000000000000001","110000001100000001",
	"110000011000000001","110000000000000010","110000001100000010","110000011000000010",
	"110000000000000011","110000001100000011","110000011000000011","110000000100000100",
	"110000001000000100","110000010000000100","110000010100000100","110000000000000000",
	"110000000000000001","110000000000000010","110000010100000010","110000011000000010",
	"110000000000000011","110000001100000011","110000010000000011","110000000000000100",
	"110000000100000100","110000001000000100","110000000100000000","110000001000000000",
	"110000001100000000","110000010000000000","110000010100000000","110000000000000001",
	"110000001100000001","110000011000000001","110000000000000010","110000001100000010",
	"110000011000000010","110000000000000011","110000001100000011","110000011000000011",
	"110000000100000100","110000010000000100","110000010100000100","110000000000000000",
	"110000000100000000","110000001000000000","110000010100000000","110000000000000001",
	"110000001000000001","110000011000000001","110000000000000010","110000001000000010",
	"110000011000000010","110000000000000011","110000001000000011","110000011000000011",
	"110000000000000100","110000001100000100","110000010000000100","110000010100000100",
	"110000001100000000","110000010000000000","110000001000000001","110000010000000001",
	"110000000100000010","110000010000000010","110000000000000011","110000000100000011",
	"110000001000000011","110000001100000011","110000010000000011","110000010100000011",
	"110000011000000011","110000010000000100","110000000100000000","110000010100000000",
	"110000000000000001","110000011000000001","110000000000000010","110000001100000010",
	"110000011000000010","110000000000000011","110000001100000011","110000011000000011",
	"110000000100000100","110000001000000100","110000010000000100","110000010100000100",
	"110000000100000000","110000011000000000","110000000000000001","110000010100000001",
	"110000011000000001","110000000000000010","110000010000000010","110000011000000010",
	"110000000000000011","110000001100000011","110000011000000011","110000000100000100",
	"110000001000000100","110000011000000100","110000000100000001","110000011000000001",
	"110000000000000010","110000000100000010","110000001000000010","110000001100000010",
	"110000010000000010","110000010100000010","110000011000000010","110000011000000011",
	"110000000100000000","110000001000000000","110000001100000000","110000010000000000",
	"110000010100000000","110000000000000001","110000011000000001","110000000000000010",
	"110000011000000010","110000000000000011","110000011000000011","110000000100000100",
	"110000001000000100","110000001100000100","110000010000000100","110000010100000100"
);
begin
	Process(CLK)
	begin
		if(CLK'event and CLK='1')then
			DATA_OUT <= M(TO_INTEGER(UNSIGNED(ADDR_OUT)));
			if(WE='1')then
				M(TO_INTEGER(UNSIGNED(ADDR_IN))) <= DATA_IN;
			end if;
		end if;
	end process;
end Behavioral;
