library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
entity ROM_DESSINS is Port (
	CLK      : in  STD_LOGIC;
	RESET    : in  STD_LOGIC;
	ADDR_OUT : in  STD_LOGIC_VECTOR (9 downto 0);
	DATA_OUT : out STD_LOGIC_VECTOR (17 downto 0);
	ADDR_IN  : in  STD_LOGIC_VECTOR (9 downto 0);
	DATA_IN  : in STD_LOGIC_VECTOR (17 downto 0);
	WE       : in  STD_LOGIC
); 
end ROM_DESSINS;
--0--\0.bmp
--1--\1.bmp
--2--\2.bmp
--3--\3.bmp
--4--\4.bmp
--5--\5.bmp
--6--\6.bmp
--7--\7.bmp
--8--\8.bmp
--9--\9.bmp
--10--\a.bmp
--11--\b.bmp
--12--\c.bmp
--13--\d.bmp
--14--\e.bmp
--15--\f.bmp
--16--\g.bmp
--17--\h.bmp
--18--\i.bmp
--19--\j.bmp
--20--\k.bmp
--21--\l.bmp
--22--\m.bmp
--23--\n.bmp
--24--\o.bmp
--25--\p.bmp
--26--\q.bmp
--27--\r.bmp
--28--\s.bmp
--29--\t.bmp
--30--\u.bmp
--31--\v.bmp
--32--\w.bmp
--33--\x.bmp
--34--\y.bmp
--35--\z.bmp
--36--\ZBALL.bmp
--37--\ZDOWN.bmp
--38--\ZLEFT.bmp
--39--\ZRIGHT.bmp
--40--\ZUP.bmp

architecture Behavioral of ROM_DESSINS is
TYPE memoire IS ARRAY(0 to 1023) OF STD_LOGIC_VECTOR(17 downto 0);--RAMBLOCK 
SIGNAL M : memoire := (
	"000100001111110000","000010101111100110","000011101111011000","000011101111001010",
	"000011101110111100","000100011110101011","000100011110011010","000010111110001111",
	"000100011101111110","000100011101101101","000100001101011101","000101001101001001",
	"000011011100111100","000100001100101100","000100011100011011","000011101100001101",
	"000100011011111100","000100011011101011","000010111011100000","000011001011010100",
	"000011111011000101","000010111010111010","000100101010101000","000101001010010100",
	"000100001010000100","000011111001110101","000100011001100100","000100101001010010",
	"000011111001000011","000010111000111000","000011111000101001","000011011000011100",
	"000100011000001011","000011010111111110","000010110111110011","000011110111100100",
	"000111000111001000","000101000110110100","000101000110100000","000101000110001100",
	"000101000101111000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"000000000000000000","000000000000000000","000000000000000000","000000000000000000",
	"111000010100000000","111000010000000001","111000001100000010","111000001000000011",
	"111000000100000100","111000000000000101","111000000100000101","111000001000000101",
	"111000001100000101","111000010000000101","111000010100000101","111000011000000101",
	"111000011100000101","111000100000000101","111000100100000101","111000000100000110",
	"111000001000000111","111000001100001000","111000010000001001","111000010100001010",
	"111000010100000000","111000010100000001","111000010100000010","111000010100000011",
	"111000000000000100","111000010100000100","111000101000000100","111000000100000101",
	"111000010100000101","111000100100000101","111000001000000110","111000010100000110",
	"111000100000000110","111000001100000111","111000010100000111","111000011100000111",
	"111000010000001000","111000010100001000","111000011000001000","111000010100001001",
	"111000010100000000","111000010000000001","111000010100000001","111000011000000001",
	"111000001100000010","111000010100000010","111000011100000010","111000001000000011",
	"111000010100000011","111000100000000011","111000000100000100","111000010100000100",
	"111000100100000100","111000000000000101","111000010100000101","111000101000000101",
	"111000010100000110","111000010100000111","111000010100001000","111000010100001001",
	"111000010000000000","111000010100000001","111000011000000010","111000011100000011",
	"111000100000000100","111000000000000101","111000000100000101","111000001000000101",
	"111000001100000101","111000010000000101","111000010100000101","111000011000000101",
	"111000011100000101","111000100000000101","111000100100000101","111000100000000110",
	"111000011100000111","111000011000001000","111000010100001001","111000010000001010",
	"111000001100000000","111000010000000000","111000010100000000","111000011000000000",
	"111000011100000000","111000001000000001","111000100000000001","111000000100000010",
	"111000100100000010","111000000000000011","111000101000000011","111000000000000100",
	"111000101000000100","111000000000000101","111000101000000101","111000000000000110",
	"111000101000000110","111000000000000111","111000101000000111","111000000100001000",
	"111000100100001000","111000001000001001","111000100000001001","111000001100001010",
	"111000010000001010","111000010100001010","111000011000001010","111000011100001010",
	"111000000000000000","111000010100000000","111000011000000000","111000000000000001",
	"111000010000000001","111000011000000001","111000000000000010","111000001100000010",
	"111000011000000010","111000000000000011","111000001000000011","111000011000000011",
	"111000000000000100","111000000100000100","111000011000000100","111000000000000000",
	"111000000100000000","111000001000000001","111000001100000001","111000010000000010",
	"111000010100000010","111000011000000010","111000001000000011","111000001100000011",
	"111000000000000100","111000000100000100","111000000000000000","111000000100000000",
	"111000010100000000","111000011000000000","111000001000000001","111000010000000001",
	"111000001100000010","111000001000000011","111000010000000011","111000000000000100",
	"111000000100000100","111000010100000100","111000011000000100","111000000000000000",
	"111000000100000000","111000001000000000","111000001100000000","111000010000000000",
	"111000010100000000","111000011000000001","111000001100000010","111000010000000010",
	"111000010100000010","111000011000000011","111000000000000100","111000000100000100",
	"111000001000000100","111000001100000100","111000010000000100","111000010100000100",
	"111000000000000000","111000000100000000","111000001000000000","111000001100000001",
	"111000010000000001","111000010100000001","111000011000000010","111000001100000011",
	"111000010000000011","111000010100000011","111000000000000100","111000000100000100",
	"111000001000000100","111000000000000000","111000000100000000","111000001000000000",
	"111000001100000000","111000010000000000","111000010100000000","111000011000000001",
	"111000011000000010","111000011000000011","111000000000000100","111000000100000100",
	"111000001000000100","111000001100000100","111000010000000100","111000010100000100",
	"111000000000000000","111000000000000001","111000000000000010","111000000100000010",
	"111000001000000010","111000001100000010","111000010000000010","111000010100000010",
	"111000011000000010","111000000000000011","111000000000000100","111000000100000000",
	"111000001000000000","111000010100000000","111000000000000001","111000001100000001",
	"111000011000000001","111000000000000010","111000001100000010","111000011000000010",
	"111000000000000011","111000001100000011","111000011000000011","111000000100000100",
	"111000010000000100","111000010100000100","111000000000000000","111000000100000000",
	"111000001000000000","111000001100000000","111000010000000000","111000010100000000",
	"111000011000000000","111000000000000001","111000001100000001","111000000000000010",
	"111000001100000010","111000010000000010","111000000000000011","111000001100000011",
	"111000010100000011","111000000100000100","111000001000000100","111000011000000100",
	"111000000100000000","111000001000000000","111000001100000000","111000010000000000",
	"111000010100000000","111000000000000001","111000011000000001","111000000000000010",
	"111000010000000010","111000011000000010","111000000000000011","111000010100000011",
	"111000000100000100","111000001000000100","111000001100000100","111000010000000100",
	"111000011000000100","111000000000000000","111000000100000000","111000001000000000",
	"111000001100000000","111000010000000000","111000010100000000","111000011000000000",
	"111000000000000001","111000001100000001","111000000000000010","111000001100000010",
	"111000000000000011","111000001100000011","111000000100000100","111000001000000100",
	"111000000100000000","111000001000000000","111000001100000000","111000010000000000",
	"111000010100000000","111000000000000001","111000011000000001","111000000000000010",
	"111000011000000010","111000000000000011","111000011000000011","111000000100000100",
	"111000001000000100","111000001100000100","111000010000000100","111000010100000100",
	"111000000000000000","111000000100000000","111000001000000000","111000001100000000",
	"111000010000000000","111000010100000000","111000011000000000","111000000100000001",
	"111000001000000001","111000001100000010","111000010000000010","111000010100000011",
	"111000011000000011","111000000000000100","111000000100000100","111000001000000100",
	"111000001100000100","111000010000000100","111000010100000100","111000011000000100",
	"111000000000000000","111000000100000000","111000001000000000","111000001100000000",
	"111000010000000000","111000010100000000","111000011000000000","111000000100000001",
	"111000001000000010","111000001100000010","111000000100000011","111000000000000100",
	"111000000100000100","111000001000000100","111000001100000100","111000010000000100",
	"111000010100000100","111000011000000100","111000000000000000","111000000100000000",
	"111000001000000000","111000001100000000","111000010000000000","111000010100000000",
	"111000011000000000","111000011000000001","111000011000000010","111000011000000011",
	"111000011000000100","111000000000000000","111000000100000000","111000001000000000",
	"111000001100000000","111000010000000000","111000010100000000","111000011000000000",
	"111000001100000001","111000001000000010","111000010000000010","111000000100000011",
	"111000010100000011","111000000000000100","111000010100000100","111000011000000100",
	"111000010000000000","111000010100000000","111000011000000001","111000011000000010",
	"111000000000000011","111000011000000011","111000000000000100","111000000100000100",
	"111000001000000100","111000001100000100","111000010000000100","111000010100000100",
	"111000000000000001","111000011000000001","111000000000000010","111000000100000010",
	"111000001000000010","111000001100000010","111000010000000010","111000010100000010",
	"111000011000000010","111000000000000011","111000011000000011","111000000000000000",
	"111000000100000000","111000001000000000","111000001100000000","111000010000000000",
	"111000010100000000","111000011000000000","111000001100000001","111000001100000010",
	"111000001100000011","111000000000000100","111000000100000100","111000001000000100",
	"111000001100000100","111000010000000100","111000010100000100","111000011000000100",
	"111000000100000000","111000001000000000","111000001100000000","111000010000000000",
	"111000010100000000","111000000000000001","111000011000000001","111000000000000010",
	"111000010000000010","111000011000000010","111000000000000011","111000010000000011",
	"111000010100000011","111000000100000100","111000010000000100","111000010100000100",
	"111000011000000100","111000000000000000","111000000100000000","111000001000000000",
	"111000001100000000","111000010000000000","111000010100000000","111000011000000000",
	"111000000000000001","111000001100000001","111000000000000010","111000001100000010",
	"111000000000000011","111000001100000011","111000000000000100","111000000000000000",
	"111000000100000000","111000001000000000","111000001100000000","111000010000000000",
	"111000010100000000","111000011000000000","111000000000000001","111000001100000001",
	"111000011000000001","111000000000000010","111000001100000010","111000011000000010",
	"111000000000000011","111000011000000011","111000000000000100","111000011000000100",
	"111000000000000000","111000000100000000","111000001000000000","111000001100000000",
	"111000010000000000","111000010100000000","111000011000000000","111000000000000001",
	"111000011000000001","111000000000000010","111000011000000010","111000000100000011",
	"111000010100000011","111000001000000100","111000001100000100","111000010000000100",
	"111000000100000000","111000001000000000","111000001100000000","111000010000000000",
	"111000010100000000","111000000000000001","111000011000000001","111000000000000010",
	"111000011000000010","111000000000000011","111000011000000011","111000000100000100",
	"111000010100000100","111000000000000000","111000000100000000","111000001000000000",
	"111000001100000000","111000010000000000","111000010100000000","111000011000000000",
	"111000000000000001","111000001100000001","111000011000000001","111000000000000010",
	"111000001100000010","111000011000000010","111000000000000011","111000001100000011",
	"111000011000000011","111000000100000100","111000001000000100","111000010000000100",
	"111000010100000100","111000001100000000","111000010000000000","111000010100000000",
	"111000011000000000","111000000100000001","111000001000000001","111000010000000001",
	"111000000000000010","111000010000000010","111000000100000011","111000001000000011",
	"111000010000000011","111000001100000100","111000010000000100","111000010100000100",
	"111000011000000100","111000000100000000","111000001000000000","111000010100000000",
	"111000000000000001","111000001100000001","111000011000000001","111000000000000010",
	"111000001100000010","111000011000000010","111000000000000011","111000001100000011",
	"111000011000000011","111000000100000100","111000001000000100","111000001100000100",
	"111000010000000100","111000010100000100","111000000100000000","111000001000000000",
	"111000010000000000","111000010100000000","111000000000000001","111000001100000001",
	"111000011000000001","111000000000000010","111000001100000010","111000011000000010",
	"111000000000000011","111000001100000011","111000011000000011","111000000100000100",
	"111000001000000100","111000010000000100","111000010100000100","111000000000000000",
	"111000000000000001","111000000000000010","111000010100000010","111000011000000010",
	"111000000000000011","111000001100000011","111000010000000011","111000000000000100",
	"111000000100000100","111000001000000100","111000000100000000","111000001000000000",
	"111000001100000000","111000010000000000","111000010100000000","111000000000000001",
	"111000001100000001","111000011000000001","111000000000000010","111000001100000010",
	"111000011000000010","111000000000000011","111000001100000011","111000011000000011",
	"111000000100000100","111000010000000100","111000010100000100","111000000000000000",
	"111000000100000000","111000001000000000","111000010100000000","111000000000000001",
	"111000001000000001","111000011000000001","111000000000000010","111000001000000010",
	"111000011000000010","111000000000000011","111000001000000011","111000011000000011",
	"111000000000000100","111000001100000100","111000010000000100","111000010100000100",
	"111000001100000000","111000010000000000","111000001000000001","111000010000000001",
	"111000000100000010","111000010000000010","111000000000000011","111000000100000011",
	"111000001000000011","111000001100000011","111000010000000011","111000010100000011",
	"111000011000000011","111000010000000100","111000000100000000","111000010100000000",
	"111000000000000001","111000011000000001","111000000000000010","111000001100000010",
	"111000011000000010","111000000000000011","111000001100000011","111000011000000011",
	"111000000100000100","111000001000000100","111000010000000100","111000010100000100",
	"111000000100000000","111000011000000000","111000000000000001","111000010100000001",
	"111000011000000001","111000000000000010","111000010000000010","111000011000000010",
	"111000000000000011","111000001100000011","111000011000000011","111000000100000100",
	"111000001000000100","111000011000000100","111000000100000001","111000011000000001",
	"111000000000000010","111000000100000010","111000001000000010","111000001100000010",
	"111000010000000010","111000010100000010","111000011000000010","111000011000000011",
	"111000000100000000","111000001000000000","111000001100000000","111000010000000000",
	"111000010100000000","111000000000000001","111000011000000001","111000000000000010",
	"111000011000000010","111000000000000011","111000011000000011","111000000100000100",
	"111000001000000100","111000001100000100","111000010000000100","111000010100000100"
);
begin
	Process(CLK)
	begin
		if(CLK'event and CLK='1')then
			DATA_OUT <= M(TO_INTEGER(UNSIGNED(ADDR_OUT)));
			if(WE='1')then
				M(TO_INTEGER(UNSIGNED(ADDR_IN))) <= DATA_IN;
			end if;
		end if;
	end process;
end Behavioral;
